module adder(a,b,c);
input [9:0]a,b;
output [9:0]c;

assign c = a + b;

endmodule
